*** SPICE deck for cell INV{lay} from library INV
*** Created on Sun Jan 26, 2014 11:32:14
*** Last revised on Sun Jan 26, 2014 12:01:48
*** Written on Sun Jan 26, 2014 12:02:40 by Electric VLSI Design System, 
*version 8.10
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
.OPTIONS NOMOD NOPAGE
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
+LVLCOD=1
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

*** TOP LEVEL CELL: INV:INV{lay}
Mnmos@2 OUT IN gnd gnd N L=0.6U W=1.5U AS=2.43P AD=3.78P PS=6.6U PD=8.1U
Mpmos@2 OUT IN vdd vdd P L=0.6U W=3U AS=5.13P AD=3.78P PS=9.6U PD=8.1U
.END
